module hw6_10();
input
output

endmodule

