module divider_tb;
parameter n = 8;
reg rem;
initial begin 
rem = 0;
