module muxdff_tb;
muxdff R0(D0, D1, Sel, Clock, Q)
endmodule